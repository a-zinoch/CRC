// 0 : CRC-32 / MPEG-2 -----------------------------------------------------------------------------
// CRC polynomial coefficients: x^32 + x^26 + x^23 + x^22 + x^16 + x^12 + x^11 + x^10 + x^8 + x^7 + x^5 + x^4 + x^2 + x + 1
//                              0x4C11DB7 (hex)
// CRC width:                   32 bits
// CRC shift direction:         left (big endian)
// Input word width:            32 bits
// ---------------------------------------------------------------------------------

// 1 : CRC-32Q ------------------------------------------------------------------------------
// CRC polynomial coefficients: x^32 + x^31 + x^24 + x^22 + x^16 + x^14 + x^8 + x^7 + x^5 + x^3 + x + 1
//                              0x814141AB (hex)
// CRC width:                   32 bits
// CRC shift direction:         left (big endian)
// Input word width:            32 bits
// ---------------------------------------------------------------------------------
module CRC32_comb(
	    input       [31:0]  data_i,
      input       [31:0]  initCrc_i,
	    input               select_i,
	    output      [31:0]  crc_o
			);

wire [31:0]CRC_0;
wire [31:0]CRC_1;

assign crc_o = select_i ? CRC_1 : CRC_0;

// CRC-32 / MPEG-2 ----------------------------------------------------------------------

assign CRC_0[0] 	= initCrc_i[0] ^ initCrc_i[6] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[12] ^ initCrc_i[16] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[12] ^ data_i[16] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31];
assign CRC_0[1] 	= initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[9] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[24] ^ initCrc_i[27] ^ initCrc_i[28] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[16] ^ data_i[17] ^ data_i[24] ^ data_i[27] ^ data_i[28];
assign CRC_0[2] 	= initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[24] ^ data_i[26] ^ data_i[30] ^ data_i[31];
assign CRC_0[3] 	= initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[25] ^ data_i[27] ^ data_i[31];
assign CRC_0[4] 	= initCrc_i[0] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[6] ^ initCrc_i[8] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[15] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[29] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[15] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[29] ^ data_i[30] ^ data_i[31];
assign CRC_0[5] 	= initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[10] ^ initCrc_i[13] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[24] ^ initCrc_i[28] ^ initCrc_i[29] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[28] ^ data_i[29];
assign CRC_0[6] 	= initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[11] ^ initCrc_i[14] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[25] ^ initCrc_i[29] ^ initCrc_i[30] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[25] ^ data_i[29] ^ data_i[30];
assign CRC_0[7] 	= initCrc_i[0] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[5] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[10] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[28] ^ initCrc_i[29] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[15] ^ data_i[16] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[28] ^ data_i[29];
assign CRC_0[8] 	= initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[8] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[17] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[28] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[17] ^ data_i[22] ^ data_i[23] ^ data_i[28] ^ data_i[31];
assign CRC_0[9] 	= initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[9] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[18] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[29] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[18] ^ data_i[23] ^ data_i[24] ^ data_i[29];
assign CRC_0[10] 	= initCrc_i[0] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[5] ^ initCrc_i[9] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[19] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[0] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[19] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_0[11] 	= initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[9] ^ initCrc_i[12] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[20] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[9] ^ data_i[12] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[20] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[31];
assign CRC_0[12] 	= initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[9] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[21] ^ initCrc_i[24] ^ initCrc_i[27] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30] ^ data_i[31];
assign CRC_0[13] 	= initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[10] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[22] ^ initCrc_i[25] ^ initCrc_i[28] ^ initCrc_i[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[22] ^ data_i[25] ^ data_i[28] ^ data_i[31];
assign CRC_0[14] 	= initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[11] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[23] ^ initCrc_i[26] ^ initCrc_i[29] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[23] ^ data_i[26] ^ data_i[29];
assign CRC_0[15] 	= initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[12] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[24] ^ initCrc_i[27] ^ initCrc_i[30] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[27] ^ data_i[30];
assign CRC_0[16] 	= initCrc_i[0] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[8] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[17] ^ initCrc_i[19] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[29] ^ initCrc_i[30] ^ data_i[0] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[12] ^ data_i[13] ^ data_i[17] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[29] ^ data_i[30];
assign CRC_0[17] 	= initCrc_i[1] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[9] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[1] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[14] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[30] ^ data_i[31];
assign CRC_0[18] 	= initCrc_i[2] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[10] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[19] ^ initCrc_i[21] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[31] ^ data_i[2] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[15] ^ data_i[19] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[28] ^ data_i[31];
assign CRC_0[19] 	= initCrc_i[3] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[11] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[29] ^ data_i[3] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[16] ^ data_i[20] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[29];
assign CRC_0[20] 	= initCrc_i[4] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[12] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[21] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[30] ^ data_i[4] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[16] ^ data_i[17] ^ data_i[21] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[30];
assign CRC_0[21] 	= initCrc_i[5] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[13] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[13] ^ data_i[17] ^ data_i[18] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
assign CRC_0[22] 	= initCrc_i[0] ^ initCrc_i[9] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[0] ^ data_i[9] ^ data_i[11] ^ data_i[12] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
assign CRC_0[23] 	= initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[6] ^ initCrc_i[9] ^ initCrc_i[13] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[6] ^ data_i[9] ^ data_i[13] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[31];
assign CRC_0[24] 	= initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[7] ^ initCrc_i[10] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[30] ^ data_i[1] ^ data_i[2] ^ data_i[7] ^ data_i[10] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[27] ^ data_i[28] ^ data_i[30];
assign CRC_0[25] 	= initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[8] ^ initCrc_i[11] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[2] ^ data_i[3] ^ data_i[8] ^ data_i[11] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_0[26] 	= initCrc_i[0] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[6] ^ initCrc_i[10] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[31] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[6] ^ data_i[10] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[31];
assign CRC_0[27] 	= initCrc_i[1] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[7] ^ initCrc_i[11] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[29];
assign CRC_0[28] 	= initCrc_i[2] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[8] ^ initCrc_i[12] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[30] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[30];
assign CRC_0[29] 	= initCrc_i[3] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[9] ^ initCrc_i[13] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[13] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_0[30] 	= initCrc_i[4] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[10] ^ initCrc_i[14] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[30] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[14] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30];
assign CRC_0[31] 	= initCrc_i[5] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[11] ^ initCrc_i[15] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[15] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[30] ^ data_i[31];

// ----------------------------------------------------------------------

// CRC-32Q ------------------------------------------------------------------ 

assign CRC_1[0]  = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[31];
assign CRC_1[1]  = initCrc_i[0] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[31] ^ data_i[0] ^ data_i[8] ^ data_i[9] ^ data_i[17] ^ data_i[18] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[31];
assign CRC_1[2]  = initCrc_i[1] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ data_i[1] ^ data_i[9] ^ data_i[10] ^ data_i[18] ^ data_i[19] ^ data_i[26] ^ data_i[27] ^ data_i[29];
assign CRC_1[3]  = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[9] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[28] ^ data_i[30] ^ data_i[31];
assign CRC_1[4]  = initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[10] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[19] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[1] ^ data_i[2] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[7] ^ data_i[8] ^ data_i[10] ^ data_i[13] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[19] ^ data_i[22] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[29] ^ data_i[31];
assign CRC_1[5]  = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[4] ^ initCrc_i[8] ^ initCrc_i[10] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[17] ^ initCrc_i[19] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[4] ^ data_i[8] ^ data_i[10] ^ data_i[12] ^ data_i[13] ^ data_i[17] ^ data_i[19] ^ data_i[21] ^ data_i[22] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[31];
assign CRC_1[6]  = initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[5] ^ initCrc_i[9] ^ initCrc_i[11] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[1] ^ data_i[2] ^ data_i[5] ^ data_i[9] ^ data_i[11] ^ data_i[13] ^ data_i[14] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[23] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_1[7]  = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[7] ^ initCrc_i[9] ^ initCrc_i[11] ^ initCrc_i[13] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[26] ^ initCrc_i[29] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[9] ^ data_i[11] ^ data_i[13] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[26] ^ data_i[29] ^ data_i[30] ^ data_i[31];
assign CRC_1[8]  = initCrc_i[0] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[11] ^ initCrc_i[13] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[30] ^ data_i[0] ^ data_i[3] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[9] ^ data_i[11] ^ data_i[13] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[30];
assign CRC_1[9]  = initCrc_i[1] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[12] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[21] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[31] ^ data_i[1] ^ data_i[4] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[12] ^ data_i[14] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[31];
assign CRC_1[10] = initCrc_i[2] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[13] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[28] ^ data_i[2] ^ data_i[5] ^ data_i[6] ^ data_i[9] ^ data_i[10] ^ data_i[11] ^ data_i[13] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[28];
assign CRC_1[11] = initCrc_i[3] ^ initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[29] ^ data_i[3] ^ data_i[6] ^ data_i[7] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[29];
assign CRC_1[12] = initCrc_i[4] ^ initCrc_i[7] ^ initCrc_i[8] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[30] ^ data_i[4] ^ data_i[7] ^ data_i[8] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[15] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[26] ^ data_i[28] ^ data_i[30];
assign CRC_1[13] = initCrc_i[5] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[5] ^ data_i[8] ^ data_i[9] ^ data_i[12] ^ data_i[13] ^ data_i[14] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[27] ^ data_i[29] ^ data_i[31];
assign CRC_1[14] = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[7] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[7] ^ data_i[11] ^ data_i[12] ^ data_i[16] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[31];
assign CRC_1[15] = initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[8] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[21] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[12] ^ data_i[13] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_1[16] = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[21] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[15] ^ data_i[16] ^ data_i[21] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[30] ^ data_i[31];
assign CRC_1[17] = initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[1] ^ data_i[2] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[16] ^ data_i[17] ^ data_i[22] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[31];
assign CRC_1[18] = initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[2] ^ data_i[3] ^ data_i[12] ^ data_i[13] ^ data_i[14] ^ data_i[17] ^ data_i[18] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_1[19] = initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[30] ^ data_i[3] ^ data_i[4] ^ data_i[13] ^ data_i[14] ^ data_i[15] ^ data_i[18] ^ data_i[19] ^ data_i[24] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[30];
assign CRC_1[20] = initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[4] ^ data_i[5] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[19] ^ data_i[20] ^ data_i[25] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[31];
assign CRC_1[21] = initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[17] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[5] ^ data_i[6] ^ data_i[15] ^ data_i[16] ^ data_i[17] ^ data_i[20] ^ data_i[21] ^ data_i[26] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_1[22] = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[29] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[9] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[19] ^ data_i[20] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[29] ^ data_i[30] ^ data_i[31];
assign CRC_1[23] = initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[14] ^ data_i[15] ^ data_i[16] ^ data_i[18] ^ data_i[20] ^ data_i[21] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[30] ^ data_i[31];
assign CRC_1[24] = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[20] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[27] ^ initCrc_i[28] ^ data_i[0] ^ data_i[1] ^ data_i[9] ^ data_i[10] ^ data_i[17] ^ data_i[18] ^ data_i[20] ^ data_i[23] ^ data_i[24] ^ data_i[25] ^ data_i[27] ^ data_i[28];
assign CRC_1[25] = initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[21] ^ initCrc_i[24] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[28] ^ initCrc_i[29] ^ data_i[1] ^ data_i[2] ^ data_i[10] ^ data_i[11] ^ data_i[18] ^ data_i[19] ^ data_i[21] ^ data_i[24] ^ data_i[25] ^ data_i[26] ^ data_i[28] ^ data_i[29];
assign CRC_1[26] = initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[22] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[29] ^ initCrc_i[30] ^ data_i[2] ^ data_i[3] ^ data_i[11] ^ data_i[12] ^ data_i[19] ^ data_i[20] ^ data_i[22] ^ data_i[25] ^ data_i[26] ^ data_i[27] ^ data_i[29] ^ data_i[30];
assign CRC_1[27] = initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[23] ^ initCrc_i[26] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[3] ^ data_i[4] ^ data_i[12] ^ data_i[13] ^ data_i[20] ^ data_i[21] ^ data_i[23] ^ data_i[26] ^ data_i[27] ^ data_i[28] ^ data_i[30] ^ data_i[31];
assign CRC_1[28] = initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[24] ^ initCrc_i[27] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[31] ^ data_i[4] ^ data_i[5] ^ data_i[13] ^ data_i[14] ^ data_i[21] ^ data_i[22] ^ data_i[24] ^ data_i[27] ^ data_i[28] ^ data_i[29] ^ data_i[31];
assign CRC_1[29] = initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[28] ^ initCrc_i[29] ^ initCrc_i[30] ^ data_i[5] ^ data_i[6] ^ data_i[14] ^ data_i[15] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[28] ^ data_i[29] ^ data_i[30];
assign CRC_1[30] = initCrc_i[6] ^ initCrc_i[7] ^ initCrc_i[15] ^ initCrc_i[16] ^ initCrc_i[23] ^ initCrc_i[24] ^ initCrc_i[26] ^ initCrc_i[29] ^ initCrc_i[30] ^ initCrc_i[31] ^ data_i[6] ^ data_i[7] ^ data_i[15] ^ data_i[16] ^ data_i[23] ^ data_i[24] ^ data_i[26] ^ data_i[29] ^ data_i[30] ^ data_i[31];
assign CRC_1[31] = initCrc_i[0] ^ initCrc_i[1] ^ initCrc_i[2] ^ initCrc_i[3] ^ initCrc_i[4] ^ initCrc_i[5] ^ initCrc_i[6] ^ initCrc_i[8] ^ initCrc_i[9] ^ initCrc_i[10] ^ initCrc_i[11] ^ initCrc_i[12] ^ initCrc_i[13] ^ initCrc_i[14] ^ initCrc_i[15] ^ initCrc_i[17] ^ initCrc_i[18] ^ initCrc_i[19] ^ initCrc_i[20] ^ initCrc_i[21] ^ initCrc_i[22] ^ initCrc_i[23] ^ initCrc_i[25] ^ initCrc_i[26] ^ initCrc_i[30] ^ data_i[0] ^ data_i[1] ^ data_i[2] ^ data_i[3] ^ data_i[4] ^ data_i[5] ^ data_i[6] ^ data_i[8] ^ data_i[9] ^ data_i[10] ^ data_i[11] ^ data_i[12] ^ data_i[13] ^ data_i[14] ^ data_i[15] ^ data_i[17] ^ data_i[18] ^ data_i[19] ^ data_i[20] ^ data_i[21] ^ data_i[22] ^ data_i[23] ^ data_i[25] ^ data_i[26] ^ data_i[30];

// ------------------------------------------------------------------------------------------

endmodule
