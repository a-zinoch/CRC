`ifndef DEFINES
`define DEFINES

	`define	PAW    				 'd8

	// CRC
  `define CRC_DATA_ADR 	 8'hD0
  `define CRC_CONF_ADR	 8'hC0
  `define CRC_OUT_ADR  	 8'hA0
  `define CRC_COUNT_ADR	 8'hA1

`endif //DEFINES